`include "kt_cache_params.sv"
`include "kt_cache.sv"
`include "sp_bram.sv"
